`timescale 1ns / 1ps
/*

    This is the module for holding the lut containing the possible duty cycle values
Unedited Table doing a whole 310Hz Sine Wave, values are split among 110 entries    
SinLut[0] = 0;
SinLut[0] =-0.0574136;
SinLut[0] =-0.114638;
SinLut[0] =-0.171484;
SinLut[0] =-0.227764;
SinLut[0] =-0.283293;
SinLut[0] =-0.337887;
SinLut[0] =-0.391367;
SinLut[0] =-0.443555;
SinLut[0] =-0.494281;
SinLut[0] =-0.543375;
SinLut[0] =-0.590677;
SinLut[0] =-0.63603;
SinLut[0] =-0.679285;
SinLut[0] =-0.720299;
SinLut[0] =-0.758937;
SinLut[0] =-0.79507;
SinLut[0] =-0.828581;
SinLut[0] =-0.859359;
SinLut[0] =-0.887301;
SinLut[0] =-0.912316;
SinLut[0] =-0.934321;
SinLut[0] =-0.953244;
SinLut[0] =-0.969022;
SinLut[0] =-0.981603;
SinLut[0] =-0.990946;
SinLut[0] =-0.99702;
SinLut[0] =-0.999804;
SinLut[0] =-0.999291;
SinLut[0] =-0.99548;
SinLut[0] =-0.988385;
SinLut[0] =-0.97803;
SinLut[0] =-0.964448;
SinLut[0] =-0.947684;
SinLut[0] =-0.927794;
SinLut[0] =-0.904843;
SinLut[0] =-0.878906;
SinLut[0] =-0.850071;
SinLut[0] =-0.81843;
SinLut[0] =-0.78409;
SinLut[0] =-0.747163;
SinLut[0] =-0.707771;
SinLut[0] =-0.666044;
SinLut[0] =-0.62212;
SinLut[0] =-0.576144;
SinLut[0] =-0.528266;
SinLut[0] =-0.478646;
SinLut[0] =-0.427447;
SinLut[0] =-0.374838;
SinLut[0] =-0.320992;
SinLut[0] =-0.266087;
SinLut[0] =-0.210304;
SinLut[0] =-0.153828;
SinLut[0] =-0.0968437;
SinLut[0] =-0.0395402;
SinLut[0] =0.0178938;
SinLut[0] =0.0752687;
SinLut[0] =0.132395;
SinLut[0] =0.189085;
SinLut[0] =0.245151;
SinLut[0] =0.300408;
SinLut[0] =0.354675;
SinLut[0] =0.407771;
SinLut[0] =0.459522;
SinLut[0] =0.509757;
SinLut[0] =0.55831;
SinLut[0] =0.605021;
SinLut[0] =0.649736;
SinLut[0] =0.692308;
SinLut[0] =0.732596;
SinLut[0] =0.770467;
SinLut[0] =0.805796;
SinLut[0] =0.838467;
SinLut[0] =0.868371;
SinLut[0] =0.895411;
SinLut[0] =0.919497;
SinLut[0] =0.940549;
SinLut[0] =0.958499;
SinLut[0] =0.973286;
SinLut[0] =0.984863;
SinLut[0] =0.99319;
SinLut[0] =0.998241;
SinLut[0] =0.999998;
SinLut[0] =0.998457;
SinLut[0] =0.993621;
SinLut[0] =0.985508;
SinLut[0] =0.974143;
SinLut[0] =0.959564;
SinLut[0] =0.94182;
SinLut[0] =0.920969;
SinLut[0] =0.897079;
SinLut[0] =0.87023;
SinLut[0] =0.84051;
SinLut[0] =0.808017;
SinLut[0] =0.772859;
SinLut[0] =0.735151;
SinLut[0] =0.695017;
SinLut[0] =0.652591;
SinLut[0] =0.608011;
SinLut[0] =0.561426;
SinLut[0] =0.512989;
SinLut[0] =0.462859;
SinLut[0] =0.411202;
SinLut[0] =0.358189;
SinLut[0] =0.303994;
SinLut[0] =0.248796;
SinLut[0] =0.192777;
SinLut[0] =0.136122;
SinLut[0] =0.0790185;
SinLut[0] =0.021654;
SinLut[0] =-0.0357819;

*/

module DutyCycle( input index,
                    output reg [0 : 31] DutyOut);
                    
reg [0 : 31] SinLut [ 0 : 120];
reg [0 : 31] counter;

initial begin
SinLut[0] = 0;
SinLut[1] =-0.0574136;
SinLut[2] =-0.114638;
SinLut[3] =-0.171484;
SinLut[4] =-0.227764;
SinLut[5] =-0.283293;
SinLut[6] =-0.337887;
SinLut[7] =-0.391367;
SinLut[8] =-0.443555;
SinLut[9] =-0.494281;
SinLut[10] =-0.543375;
SinLut[11] =-0.590677;
SinLut[12] =-0.63603;
SinLut[13] =-0.679285;
SinLut[14] =-0.720299;
SinLut[15] =-0.758937;
SinLut[16] =-0.79507;
SinLut[17] =-0.828581;
SinLut[18] =-0.859359;
SinLut[19] =-0.887301;
SinLut[20] =-0.912316;
SinLut[21] =-0.934321;
SinLut[22] =-0.969022;
SinLut[23] =-0.981603;
SinLut[24] =-0.99702;
SinLut[25] =-0.999804;
SinLut[26] =-0.999291;
SinLut[27] =-0.988385;
SinLut[28] =-0.97803;
SinLut[29] =-0.964448;
SinLut[30] =-0.947684;
SinLut[31] =-0.927794;
SinLut[32] =-0.904843;
SinLut[33] =-0.878906;
SinLut[34] =-0.850071;
SinLut[35] =-0.81843;
SinLut[36] =-0.78409;
SinLut[37] =-0.747163;
SinLut[38] =-0.707771;
SinLut[39] =-0.666044;
SinLut[40] =-0.62212;
SinLut[41] =-0.576144;
SinLut[42] =-0.528266;
SinLut[43] =-0.478646;
SinLut[44] =-0.427447;
SinLut[45] =-0.374838;
SinLut[46] =-0.320992;
SinLut[47] =-0.266087;
SinLut[48] =-0.210304;
SinLut[49] =-0.153828;
SinLut[50] =-0.0968437;
SinLut[51] =-0.0395402;
SinLut[52] =0.0178938;
SinLut[53] =0.0752687;
SinLut[54] =0.132395;
SinLut[55] =0.189085;
SinLut[56] =0.245151;
SinLut[57] =0.300408;
SinLut[58] =0.354675;
SinLut[59] =0.407771;
SinLut[60] =0.459522;
SinLut[61] =0.509757;
SinLut[62] =0.55831;
SinLut[63] =0.605021;
SinLut[64] =0.649736;
SinLut[65] =0.692308;
SinLut[66] =0.732596;
SinLut[67] =0.770467;
SinLut[68] =0.805796;
SinLut[69] =0.838467;
SinLut[70] =0.895411;
SinLut[71] =0.919497;
SinLut[72] =0.940549;
SinLut[73] =0.973286;
SinLut[74] =0.998241;
SinLut[75] =0.999998;
SinLut[76] =0.998457;
SinLut[78] =0.985508;
SinLut[79] =0.974143;
SinLut[80] =0.959564;
SinLut[81] =0.920969;
SinLut[82] =0.897079;
SinLut[83] =0.84051;
SinLut[84] =0.808017;
SinLut[85] =0.772859;
SinLut[86] =0.735151;
SinLut[87] =0.695017;
SinLut[88] =0.652591;
SinLut[89] =0.608011;
SinLut[90] =0.561426;
SinLut[91] =0.512989;
SinLut[92] =0.462859;
SinLut[93] =0.411202;
SinLut[94] =0.358189;
SinLut[95] =0.303994;
SinLut[96] =0.248796;
SinLut[97] =0.192777;
SinLut[98] =0.136122;
SinLut[99] =0.0790185;
SinLut[100] =0.021654;
SinLut[101] =0;
counter = 32'b0;
end

always @(negedge index) begin
  
   if(counter == 32'd101) begin
    counter = 32'd0;
   end
   else begin
    counter = counter + 32'd1;
   end
    DutyOut = SinLut[counter];
end

endmodule
